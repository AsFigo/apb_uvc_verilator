`define AF_NO_UVM_RAL
/* verilator lint_off REDEFMACRO */
`define uvm_field_enum(T,ARG,FLAG=UVM_DEFAULT) \
  // Dummy macro
